library verilog;
use verilog.vl_types.all;
entity contador_temp_vlg_vec_tst is
end contador_temp_vlg_vec_tst;
