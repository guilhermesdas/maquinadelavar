library verilog;
use verilog.vl_types.all;
entity ligadesliga_vlg_sample_tst is
    port(
        botao           : in     vl_logic;
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ligadesliga_vlg_sample_tst;
