library verilog;
use verilog.vl_types.all;
entity historia4_vlg_check_tst is
    port(
        off             : in     vl_logic;
        rst             : in     vl_logic;
        Standby         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end historia4_vlg_check_tst;
