library verilog;
use verilog.vl_types.all;
entity contador_divfreq_vlg_vec_tst is
end contador_divfreq_vlg_vec_tst;
