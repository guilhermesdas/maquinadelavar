library verilog;
use verilog.vl_types.all;
entity cont_divfreq_vlg_vec_tst is
end cont_divfreq_vlg_vec_tst;
