library verilog;
use verilog.vl_types.all;
entity historia2_vlg_vec_tst is
end historia2_vlg_vec_tst;
