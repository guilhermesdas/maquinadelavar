library verilog;
use verilog.vl_types.all;
entity debounce_vlg_vec_tst is
end debounce_vlg_vec_tst;
