library verilog;
use verilog.vl_types.all;
entity COMPLETA_vlg_vec_tst is
end COMPLETA_vlg_vec_tst;
