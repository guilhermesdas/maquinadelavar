library verilog;
use verilog.vl_types.all;
entity divfreq_vlg_vec_tst is
end divfreq_vlg_vec_tst;
