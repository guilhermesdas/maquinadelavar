library verilog;
use verilog.vl_types.all;
entity ligadesliga_vlg_vec_tst is
end ligadesliga_vlg_vec_tst;
