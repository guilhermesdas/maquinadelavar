library verilog;
use verilog.vl_types.all;
entity historia4_vlg_vec_tst is
end historia4_vlg_vec_tst;
